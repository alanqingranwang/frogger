module font_rom ( input [4:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 5;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x01
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
		  
        16'b0001001111001000, // 4
        16'b0011011111101100, // 5
        16'b0001011111101000, // 6
        16'b0001111111111000, // 7
        16'b0000011111100000, // 8
        16'b0001111111111000, // 9
        16'b0001011111101000, // a
        16'b0011001111001100, // b
        16'b0001000000001000, // c
		  
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
        
         // code x23
        
        };
		  
		  /*
		  16'b0001002122001000, // 4
        16'b0011031221301100, // 5
        16'b0001011221101000, // 6
        16'b0001122222211000, // 7
        16'b0000021222200000, // 8
        16'b0001121222211000, // 9
        16'b0001012122101000, // a
        16'b0011001221001100, // b
        16'b0001000000001000, // c
		  */

	assign data = ROM[addr];

endmodule 