module Sprites (  output logic [0:15][0:15][0:1]  FrogSprite,
						output logic [0:15][0:31][0:1]  TruckSprite,
						output logic [0:15][0:15][0:1]  YellowCarSprite,
						output logic [0:15][0:15][0:1]  GrayCarSprite,
						output logic [0:15][0:15][0:1]  TractorSprite,
						output logic [0:15][0:47][0:1]  FishThreeSprite,
						output logic [0:15][0:47][0:1]  LogSprite,
						output logic [0:15][0:31][0:1]  FishTwoSprite,
						output logic [0:15][0:63][0:1]  BigLogSprite,
						output logic [0:17][0:17][0:1]  SafeFrogSprite,
						output logic [0:16][0:111][0:1] TitleSprite,
						output logic [0:15][0:15][0:1]  DeathSprite,
						output logic [0:9][0:103][0:1]  Player1Sprite,
						output logic [0:9][0:103][0:1]  Player2Sprite,
						output logic [0:9][0:55][0:1]   WinSprite,
						output logic [0:9][0:71][0:1]   GameOverSprite,
						output logic [0:9][0:87][0:1]   PressEnterSprite
);

always_comb
begin

FrogSprite <= '{
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,1,0,0,2,1,2,2,0,0,1,0,0,0},
				  '{0,0,1,1,0,3,1,2,2,1,3,0,1,1,0,0},
				  '{0,0,0,1,0,1,1,2,2,1,1,0,1,0,0,0},
				  '{0,0,0,1,1,2,2,2,2,2,2,1,1,0,0,0},
				  '{0,0,0,0,0,2,1,2,2,2,2,0,0,0,0,0},
				  '{0,0,0,1,1,2,1,2,2,2,2,1,1,0,0,0},
				  '{0,0,0,1,0,1,2,1,2,2,1,0,1,0,0,0},
				  '{0,0,1,1,0,0,1,2,2,1,0,0,1,1,0,0},
				  '{0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
			};
			
TruckSprite <= '{
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},	
					'{0,0,0,0,0,3,3,3,0,0,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0},
					'{0,0,0,2,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,2,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,2,1,1,1,1,1,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,2,1,1,1,1,1,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,2,1,1,1,1,1,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,2,1,1,1,1,1,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,2,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,0,2,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					'{0,0,0,0,0,3,3,3,0,0,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
			};

YellowCarSprite <= '{
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1},
				  '{0,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1},
				  '{0,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1},
				  '{0,0,0,0,0,3,0,0,0,0,0,0,0,3,0,0},
				  '{0,0,0,2,2,2,2,2,2,2,2,2,2,2,2,0},
				  '{3,0,2,2,2,2,3,3,3,2,2,3,3,3,3,3},
				  '{0,2,2,2,2,3,3,3,2,2,1,2,1,2,1,2},
				  '{0,2,2,2,2,3,3,3,2,2,1,2,1,2,1,2},
				  '{3,0,2,2,2,2,3,3,3,2,2,3,3,3,3,3},
				  '{0,0,0,2,2,2,2,2,2,2,2,2,2,2,2,0},
				  '{0,0,0,0,0,3,0,0,0,0,0,0,0,3,0,0},
				  '{0,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1},
				  '{0,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1},
				  '{0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
				};
				
GrayCarSprite <= '{
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0},
				  '{0,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0},
				  '{0,0,3,0,0,0,0,0,0,0,0,3,0,0,0,0},
				  '{0,2,2,2,2,2,2,2,2,2,2,2,2,0,0,0},				  
				  '{0,3,3,3,3,2,2,3,3,3,2,2,2,2,0,3},
				  '{0,1,2,1,2,1,2,2,3,3,3,2,2,2,2,0},
				  '{0,1,2,1,2,1,2,2,3,3,3,2,2,2,2,0},				  
				  '{0,3,3,3,3,2,2,3,3,3,2,2,2,2,0,3},
				  '{0,2,2,2,2,2,2,2,2,2,2,2,2,0,0,0},
				  '{0,0,3,0,0,0,0,0,0,0,3,0,0,0,0,0},
				  '{0,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0},
				  '{0,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0},
				  '{0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0},
				  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
				};
				
TractorSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,3,1,3,1,3,1,3,0,0,0,0,1,1,1,0},
					  '{0,3,1,3,1,3,1,3,0,0,0,0,1,3,0,0},
					  '{0,0,2,0,0,0,2,0,0,2,2,2,1,1,1,0},
					  '{0,0,1,1,1,1,1,1,1,1,0,0,1,3,0,0},
					  '{0,1,1,1,1,1,2,2,1,2,0,0,1,1,1,0}, 
					  '{0,1,1,2,2,2,1,2,1,1,0,0,1,3,0,0},
					  '{0,1,1,2,2,2,1,2,1,1,0,0,1,3,0,0},
					  '{0,1,1,1,1,1,2,2,1,2,0,0,1,1,1,0},
					  '{0,0,1,1,1,1,1,1,1,1,0,0,1,3,0,0},
					  '{0,0,2,0,0,0,2,0,0,2,2,2,1,1,1,0},
					  '{0,1,3,1,3,1,3,1,0,0,0,0,1,3,0,0},
					  '{0,1,3,1,3,1,3,1,0,0,0,0,1,1,1,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}					  
};

FishThreeSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0},
					  '{0,0,0,2,2,3,3,3,3,3,2,2,0,0,0,0,0,0,0,2,2,3,3,3,3,3,2,2,0,0,0,0,0,0,0,2,2,3,3,3,3,3,2,2,0,0,0,0},  
					  '{0,0,0,0,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,0,0,0,0,0},		  
					  '{0,0,1,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,1,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,1,3,3,3,3,3,3,3,3,3,0,0,0,0},  
					  '{0,2,2,3,3,3,3,3,3,3,3,3,3,2,0,0,0,2,2,3,3,3,3,3,3,3,3,3,3,2,0,0,0,2,2,3,3,3,3,3,3,3,3,3,3,2,0,0}, 		  
					  '{0,0,1,3,3,3,3,3,3,3,1,3,0,0,0,0,0,0,1,3,3,3,3,3,3,3,1,3,0,0,0,0,0,0,1,3,3,3,3,3,3,3,1,3,0,0,0,0},
					  '{0,0,0,0,3,1,3,3,3,1,3,0,0,0,0,0,0,0,0,0,3,1,3,3,3,1,3,0,0,0,0,0,0,0,0,0,3,1,3,3,3,1,3,0,0,0,0,0},
					  '{0,0,0,2,2,3,1,1,1,3,2,2,0,0,0,0,0,0,0,2,2,3,1,1,1,3,2,2,0,0,0,0,0,0,0,2,2,3,1,1,1,3,2,2,0,0,0,0},		  
					  '{0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0},		  
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},					  
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}					  
					  };
					  
FishTwoSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0},
					  '{0,0,0,2,2,3,3,3,3,3,2,2,0,0,0,0,0,0,0,2,2,3,3,3,3,3,2,2,0,0,0,0},  
					  '{0,0,0,0,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,0,0,0,0,0},		  
					  '{0,0,1,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,1,3,3,3,3,3,3,3,3,3,0,0,0,0},  
					  '{0,2,2,3,3,3,3,3,3,3,3,3,3,2,0,0,0,2,2,3,3,3,3,3,3,3,3,3,3,2,0,0}, 		  
					  '{0,0,1,3,3,3,3,3,3,3,1,3,0,0,0,0,0,0,1,3,3,3,3,3,3,3,1,3,0,0,0,0},
					  '{0,0,0,0,3,1,3,3,3,1,3,0,0,0,0,0,0,0,0,0,3,1,3,3,3,1,3,0,0,0,0,0},
					  '{0,0,0,2,2,3,1,1,1,3,2,2,0,0,0,0,0,0,0,2,2,3,1,1,1,3,2,2,0,0,0,0},		  
					  '{0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0,0,0},		  
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},					  
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}					  
					  };
					  
LogSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,1,1,1,1,1,1,1,0,1,1,1,1,0,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,3,3,3,0,0,0,0,0},
					  '{0,0,0,0,1,1,1,1,1,1,3,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,3,3,3,3,3,0,0,0,0},
					  '{0,0,0,0,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,3,0,0,0,0},  
					  '{0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,3,1,1,1,3,3,0,0,0},		  
					  '{0,0,0,1,1,1,1,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1,3,0,0,0},  
					  '{0,0,0,1,1,3,3,1,1,1,1,3,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,3,1,1,3,0,0,0}, 		  
					  '{0,0,0,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,3,1,1,1,1,1,3,3,1,3,3,3,1,3,1,3,3,0,0,0},
					  '{0,0,0,0,1,1,1,1,1,1,1,0,2,3,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,2,2,2,2,2,2,2,2,3,1,1,1,3,0,0,0,0},
					  '{0,0,0,0,0,0,2,0,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,1,1,3,3,0,0,0,0},		  
					  '{0,0,0,0,0,1,1,1,2,2,2,0,2,2,2,2,2,2,2,0,2,2,2,2,2,2,2,0,2,2,2,2,2,2,2,2,0,2,2,2,1,3,3,0,0,0,0,0},		  
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
					  };
					  
BigLogSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,1,1,1,1,1,1,1,0,1,1,1,1,0,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,0,1,1,1,1,1,3,3,3,0,0,0,0,0},
					  '{0,0,0,0,1,1,1,1,1,1,3,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,3,3,3,3,3,0,0,0,0},
					  '{0,0,0,0,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,3,0,0,0,0},  
					  '{0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,3,1,1,1,3,3,0,0,0},		  
					  '{0,0,0,1,1,1,1,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1,3,0,0,0},  
					  '{0,0,0,1,1,3,3,1,1,1,1,3,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,3,1,1,3,0,0,0}, 		  
					  '{0,0,0,1,1,1,1,1,1,1,1,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,3,1,1,1,1,1,3,3,1,3,3,3,1,3,1,3,3,0,0,0},
					  '{0,0,0,0,1,1,1,1,1,1,1,0,2,3,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,2,2,2,2,2,2,2,2,3,1,1,1,3,0,0,0,0},
					  '{0,0,0,0,0,0,2,0,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,1,1,3,3,0,0,0,0},		  
					  '{0,0,0,0,0,1,1,1,2,2,2,0,2,2,2,2,2,2,2,0,2,2,2,2,2,2,2,0,2,2,2,2,2,2,2,0,2,2,2,2,2,2,2,0,2,2,2,2,2,2,2,2,0,2,2,2,1,3,3,0,0,0,0,0},		  
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
					  };
					  
SafeFrogSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,0},
					  '{0,0,0,1,0,0,1,0,0,0,0,1,0,0,1,0,0,0},
					  '{0,0,0,1,2,2,1,1,1,1,1,1,2,2,1,0,0,0},
					  '{0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0}, 
					  '{0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0},
					  '{0,0,0,0,0,1,1,2,1,1,2,1,1,0,0,0,0,0},	  
					  '{0,0,1,0,0,1,1,1,2,2,1,1,1,0,0,1,0,0},   
					  '{0,1,1,1,0,3,1,1,1,1,1,1,3,0,1,1,1,0},		  
					  '{0,1,1,1,1,3,1,1,1,1,1,1,3,1,1,1,1,0},	  
					  '{0,1,1,1,1,3,3,1,1,1,1,3,3,1,1,1,1,0},	  
					  '{0,1,1,1,1,1,3,3,3,3,3,3,1,1,1,1,1,0},
					  '{0,0,1,1,1,1,3,2,2,2,3,3,1,1,1,1,0,0},	  
					  '{0,0,1,1,1,1,3,2,2,2,3,3,1,1,1,1,0,0},		  
					  '{0,0,0,0,1,1,1,3,3,3,3,1,1,1,0,0,0,0},		  
					  '{0,0,0,1,1,1,1,0,0,0,0,1,1,1,1,0,0,0},
					  '{0,0,1,1,1,0,1,0,0,0,0,1,0,1,1,1,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};					  


TitleSprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},					  
					  '{0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					  '{0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0},
					  '{0,2,1,1,1,1,3,3,3,3,3,3,3,3,3,0,0,2,1,1,1,1,3,3,3,3,3,2,1,1,1,1,0,0,1,1,1,1,3,3,3,3,3,2,1,1,1,1,0,0,0,0,1,1,1,1,3,3,3,3,3,3,3,0,0,0,0,0,1,1,1,1,3,3,3,3,3,3,3,0,0,0,2,1,1,1,1,3,3,3,3,3,3,3,0,0,2,1,1,1,1,3,3,3,3,3,2,1,1,1,1,0},			  
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0}, 			  
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,0,1,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0},
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0},	   
					  '{0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,0,1,1,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,1,1,1,1,1,1,0,2,1,1,1,1,0,0,0,0,1,1,1,1,1,1,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,0,1,1,1,1,1,1,0},   
					  '{0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,2,1,1,1,1,1,1,0,2,1,1,1,1,0,0,0,2,1,1,1,1,1,1,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,1,1,0},				  
					  '{0,2,1,1,1,1,3,3,3,3,3,3,3,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,3,3,3,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,3,3,2,1,1,1,1,0,2,1,1,1,1,0,0,0,3,3,2,1,1,1,1,0,0,2,1,1,1,1,3,3,3,3,3,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,3,3,3,0,0},	
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0},	
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,3,3,2,1,1,1,1,0,0,0,2,1,1,1,1,0,3,3,2,1,1,1,1,0,0,0,2,1,1,1,1,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,0,0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0},			  
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,3,3,3,2,1,1,1,1,1,1,0,3,3,2,1,1,1,1,1,1,1,1,1,1,3,0,0,0,0,3,3,2,1,1,1,1,1,1,1,1,1,1,0,0,0,3,3,2,1,1,1,1,1,1,1,1,1,1,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,2,1,1,1,1,3,3,3,2,1,1,1,1,1,1,0},
					  '{0,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,2,1,1,1,1,0,0,0,2,1,1,1,1,1,1,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,2,1,1,1,1,1,1,1,1,1,1,0,0,2,1,1,1,1,1,1,1,1,1,1,1,1,0,2,1,1,1,1,0,0,0,2,1,1,1,1,1,1,0},
					  '{0,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,0,0,0,0,3,3,3,3,3,3,0,0,0,0,3,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,0,0,3,3,3,3,3,3,3,3,3,3,0,0,0,0,0,0,3,3,3,3,3,3,3,3,3,3,0,0,0,3,3,3,3,3,3,3,3,3,3,3,3,0,0,3,3,3,3,0,0,0,0,3,3,3,3,3,3,0,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}					  
};					  

DeathSprite <= '{
					  '{0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0},
					  '{0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0},
					  '{0,0,0,0,1,1,0,1,1,1,0,1,1,0,0,0},
					  '{0,0,0,0,1,0,1,1,1,1,1,0,1,0,0,0},	  
					  '{0,1,1,0,1,1,1,1,1,1,1,1,1,0,1,1}, 
					  '{0,1,1,0,0,0,1,1,1,1,1,0,0,0,1,1},	  
					  '{0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0},   	  
					  '{0,0,0,1,0,0,0,1,1,1,0,0,0,1,0,0},		  
					  '{0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0},		  
					  '{0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0},	    
					  '{0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0},  
					  '{0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0},	 
					  '{0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0},		
					  '{0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0},		  
					  '{0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0},
					  '{0,0,0,0,1,1,0,0,0,0,0,1,1,0,0,0}					  
};				

Player1Sprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,1,1,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,1,1,1,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0},
					  '{0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,1,1,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,1,1,0,0,1,1,1,0,1,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,1,1,0,0,1,1,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,1,1,0,0,1,1,0,0,0,0,0,0,1,1,0,0,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,1,0,1,1,0,1,1,1,1,1,0,0,0},
					  '{0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0,1,1,0,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,1,1,1,1,1,0,1,1,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}

};	

Player2Sprite <= '{
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
					  '{0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0, 1,1,1,1,1,1,0,0, 1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,1,1,0,0,1,1,0, 1,1,1,1,1,1,1,0, 1,1,1,1,1,1,0,0, 0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,1,1,1,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0},
					  '{1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0, 1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,1,1,0, 1,1,0,0,0,0,0,0, 1,1,0,0,0,1,1,0, 0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,1,1,0,0,1,1,1,0,1,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0, 1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,1,1,0,0,1,1,0, 1,1,0,0,0,0,0,0, 1,1,0,0,0,1,1,0, 0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0, 1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,1,1,0,0, 1,1,0,0,0,0,0,0, 1,1,0,0,1,1,1,0, 0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,0,0,0},
					  '{0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0, 1,1,1,1,1,1,0,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0, 1,1,1,1,1,0,0,0, 1,1,1,1,1,0,0,0, 0,0,0,0,0,0,0,0,1,1,0,0,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,1,0,1,1,0,1,1,1,1,1,0,0,0},
					  '{0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0, 1,1,0,0,0,0,0,0, 1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,1,1,0,0,0, 1,1,0,0,0,0,0,0, 1,1,0,1,1,1,0,0, 0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0},
					  '{1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0, 1,1,0,0,0,0,0,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0, 1,1,0,0,0,0,0,0, 1,1,0,0,1,1,1,0, 0,0,0,0,0,0,0,0,0,1,1,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0},
					  '{1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0, 1,1,0,0,0,0,0,0, 1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0, 1,1,1,1,1,1,1,0, 1,1,0,0,1,1,1,0, 0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0},
					  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}

};  

WinSprite <= '{
				 '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
				 '{0,1,1,0,0,1,1,0,0,1,1,1,1,1,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0},
				 '{0,1,1,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,1,0,0,1,1,0},
				 '{0,1,1,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,1,0,1,1,0,0,0,0,1,1,0,0,0,1,1,1,1,0,1,1,0},
				 '{0,0,1,1,1,1,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,1,1,0,0,0,1,1,1,1,1,1,1,0},
				 '{0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,1,0},
				 '{0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,1,1,1,0},
				 '{0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,1,1,0},
				 '{0,0,0,1,1,0,0,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0},
				 '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};

GameOverSprite <= '{
					   '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0},
						'{0,0,1,1,1,1,1,0,0,0,1,1,1,0,0,0,1,1,0,0,0,1,1,0, 1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0, 1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0, 1,1,1,1,1,1,0,0},
						'{0,1,1,0,0,0,0,0,0,1,1,0,1,1,0,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0, 1,1,0,0,0,1,1,0},
						'{1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,0, 1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0, 1,1,0,0,0,1,1,0},
						'{1,1,0,0,1,1,1,0,1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0, 1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,1,1,0,1,1,0,0,0,0,0,0, 1,1,0,0,1,1,1,0},
						'{1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,1,0,1,1,0, 1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0, 1,1,1,0,1,1,1,0,1,1,1,1,1,0,0,0, 1,1,1,1,1,0,0,0},
						'{1,1,0,0,0,1,1,0,1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0, 0,1,1,1,1,1,0,0,1,1,0,0,0,0,0,0, 1,1,0,1,1,1,0,0},
						'{0,1,1,0,0,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,0, 0,0,1,1,1,0,0,0,1,1,0,0,0,0,0,0, 1,1,0,0,1,1,1,0},
						'{0,0,1,1,1,1,1,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0, 1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0, 0,0,0,1,0,0,0,0,1,1,1,1,1,1,1,0, 1,1,0,0,1,1,1,0},
						'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0}

};

PressEnterSprite <= '{
						  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0},
						  '{1,1,1,1,1,1,0,0,1,1,1,1,1,1,0,0, 1,1,1,1,1,1,1,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0,0,1,1,1,1,1,1,0,1,1,1,1,1,1,1,0, 1,1,1,1,1,1,0,0},
						  '{1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,1,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0, 1,1,0,0,0,1,1,0},
						  '{1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,1,1,0,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0, 1,1,0,0,0,1,1,0},
						  '{1,1,0,0,0,1,1,0,1,1,0,0,1,1,1,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0, 1,1,0,0,1,1,1,0},
						  '{1,1,1,1,1,1,0,0,1,1,1,1,1,0,0,0, 1,1,1,1,1,0,0,0,0,1,1,1,1,1,1,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,1,1,0,1,1,1,1,0,0,0,0,1,1,0,0,0,1,1,1,1,1,0,0,0, 1,1,1,1,1,0,0,0},
						  '{1,1,0,0,0,0,0,0,1,1,0,1,1,1,0,0, 1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,1,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0, 1,1,0,1,1,1,0,0},
						  '{1,1,0,0,0,0,0,0,1,1,0,0,1,1,1,0, 1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,0,0,0,0,0,0, 1,1,0,0,1,1,1,0},
						  '{1,1,0,0,0,0,0,0,1,1,0,0,1,1,1,0, 1,1,1,1,1,1,1,0,0,1,1,1,1,1,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,1,1,0,0,0,1,1,0,0,0,0,1,1,0,0,0,1,1,1,1,1,1,1,0, 1,1,0,0,1,1,1,0},
						  '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0, 0,0,0,0,0,0,0,0}
							};


end 
endmodule
